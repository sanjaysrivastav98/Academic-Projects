module FADDER_1_beh(A,B,M,S,C);
	input A;
	input B;
	input M;
	output S;
	output C;
	
	