`include "FADDER_1.v"

module FADDER_4_beh(A,B,C,S);