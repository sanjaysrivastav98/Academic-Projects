module mux4_1(regData,q1,q2,q3,q4,reg_no);